	component accel is
		port (
			accelerometer_spi_external_interface_I2C_SDAT      : inout std_logic                    := 'X'; -- I2C_SDAT
			accelerometer_spi_external_interface_I2C_SCLK      : out   std_logic;                           -- I2C_SCLK
			accelerometer_spi_external_interface_G_SENSOR_CS_N : out   std_logic;                           -- G_SENSOR_CS_N
			accelerometer_spi_external_interface_G_SENSOR_INT  : in    std_logic                    := 'X'; -- G_SENSOR_INT
			clk_clk                                            : in    std_logic                    := 'X'; -- clk
			hex_0_export                                       : out   std_logic_vector(6 downto 0);        -- export
			hex_1_export                                       : out   std_logic_vector(6 downto 0);        -- export
			hex_2_export                                       : out   std_logic_vector(6 downto 0);        -- export
			hex_3_export                                       : out   std_logic_vector(6 downto 0);        -- export
			hex_4_export                                       : out   std_logic_vector(6 downto 0);        -- export
			hex_5_export                                       : out   std_logic_vector(6 downto 0);        -- export
			led_external_connection_export                     : out   std_logic_vector(9 downto 0);        -- export
			reset_reset_n                                      : in    std_logic                    := 'X'  -- reset_n
		);
	end component accel;

	u0 : component accel
		port map (
			accelerometer_spi_external_interface_I2C_SDAT      => CONNECTED_TO_accelerometer_spi_external_interface_I2C_SDAT,      -- accelerometer_spi_external_interface.I2C_SDAT
			accelerometer_spi_external_interface_I2C_SCLK      => CONNECTED_TO_accelerometer_spi_external_interface_I2C_SCLK,      --                                     .I2C_SCLK
			accelerometer_spi_external_interface_G_SENSOR_CS_N => CONNECTED_TO_accelerometer_spi_external_interface_G_SENSOR_CS_N, --                                     .G_SENSOR_CS_N
			accelerometer_spi_external_interface_G_SENSOR_INT  => CONNECTED_TO_accelerometer_spi_external_interface_G_SENSOR_INT,  --                                     .G_SENSOR_INT
			clk_clk                                            => CONNECTED_TO_clk_clk,                                            --                                  clk.clk
			hex_0_export                                       => CONNECTED_TO_hex_0_export,                                       --                                hex_0.export
			hex_1_export                                       => CONNECTED_TO_hex_1_export,                                       --                                hex_1.export
			hex_2_export                                       => CONNECTED_TO_hex_2_export,                                       --                                hex_2.export
			hex_3_export                                       => CONNECTED_TO_hex_3_export,                                       --                                hex_3.export
			hex_4_export                                       => CONNECTED_TO_hex_4_export,                                       --                                hex_4.export
			hex_5_export                                       => CONNECTED_TO_hex_5_export,                                       --                                hex_5.export
			led_external_connection_export                     => CONNECTED_TO_led_external_connection_export,                     --              led_external_connection.export
			reset_reset_n                                      => CONNECTED_TO_reset_reset_n                                       --                                reset.reset_n
		);

